// DMA Transaction class

typedef enum {STIMULUS,BASE_ADDR_CFG,BASE_COUNT_CFG,REG_WRITE_CFG,REG_READ_CFG} pkt_type_t;

class dma_transaction;

import dma_reg_pkg::*;

   pkt_type_t tx_type;
   
  // Properties
  // declare all inputs and controls signals as rand to generate random values from them
  rand bit ior;
  rand bit iow;
  bit [7:0] data;
  //rand bit [7:0] data_out;
  bit [3:0] addr_lo;
  //rand bit [3:0] out_addr;
  rand bit eop;
  rand bit [3:0] dreq;
  bit [3:0] dreq_old;
  bit [3:0] dack_sampled;
  rand bit hlda;
  rand bit cs;
  
 // outputs will be generated by the DUT hence no rand
  bit [3:0] addr_hi;
  bit [3:0] dack;
  bit hrq;
  bit aen;
  bit adstb;
  
  //control register write done flag
  bit ctrl_regs_wr_done;
  
  // Methods
  // deep copy method
  function void copy(output dma_transaction tx);
    tx = new;
    tx.ior = this.ior;
    tx.iow = this.iow;
    tx.data = this.data;
    tx.addr_lo = this.addr_lo;
    tx.eop = this.eop;
    tx.dreq = this.dreq;
    tx.hlda = this.hlda;
    tx.cs = this.cs;
    tx.addr_hi = this.addr_hi;
    tx.dack = this.dack;
    tx.hrq = this.hrq;
    tx.aen = this.aen;
    tx.adstb = this.adstb;
  endfunction
  
  function void compare(input dma_transaction tx);
    if(
      tx.ior != this.ior ||
      tx.iow != this.iow ||
      tx.data != this.data ||
      tx.addr_lo != this.addr_lo ||
      tx.eop != this.eop ||
      tx.dreq != this.dreq ||
      tx.hlda != this.hlda ||
      tx.cs != this.cs ||
      tx.addr_hi != this.addr_hi ||
      tx.dack != this.dack ||
      tx.hrq != this.hrq ||
      tx.aen != this.aen ||
      tx.adstb != this.adstb)
        return 0;         // compare failed
    else
        return 1;         // compare passed
  endfunction
  
  function void print();
      	$display("-----PRINTING TRANSACTION CLASS PROPERTIES---------");
      	$display("\t IOR = %b", tx.ior);
      	$display("\t IOW = %b", tx.iow);
		$display("\t DATA = %b", tx.data);
		$display("\t ADDR_L = %b", tx.addr_lo);
		$display("\t ADDR_H = %b", tx.addr_hi);
		$display("\t EOP = %b", tx.eop);
		$display("\t DREQ = %b", tx.dreq);
		$display("\t DACK = %b", tx.dack);
		$display("\t HLDA = %b", tx.hlda);
		$display("\t HRQ = %b", tx.hrq);
		$display("\t CS = %b", tx.cs);
		$display("\t AEN = %b", tx.aen);
		$display("\t ADSTB = %b", tx.adstb);
		$display("---------------------------------------------------");
  endfunction

// Initialize the registers	
task regs_init();	
	CMD_REG					= '0;
	REQ_REG					= '0;
	MASK_REG				= '0;
	STATUS_REG				= '0;
	TEMP_DATA_REG			= '0;
	foreach(MODE_REG[i])				MODE_REG[i] 			= '0;
	foreach(TEMP_ADDR_REG[i])			TEMP_ADDR_REG[i]		= '0;
	foreach(TEMP_WORD_COUNT_REG[i]) 	TEMP_WORD_COUNT_REG[i]  = '0;
	foreach(BASE_ADDR_REG[i])			BASE_ADDR_REG[i]		= '0;
	foreach(BASE_WORD_COUNT_REG[i]) 	BASE_WORD_COUNT_REG		= '0;
	foreach(CURR_ADDR_REG[i])			CURR_ADDR_REG 			= '0;
	foreach(CURR_WORD_COUNT_REG[i])		CURR_WORD_COUNT_REG		= '0;
endtask : regs_init

// TODO : confirm prototype
// Read Register
/*
task regs_read(bit[3:0] address, bit [15:0] data);
	tx = new();
	tx.pkt_type = REG_READ;
	tx.cs = 1'b0;
	tx.ior = 1'b0;
	tx.iow = 1'b1;
	tx.addr_lo = address;
	tx.dreq = 4'b0;
	tx.hlda = 1'b0;
	tx.eop = 1'b1;
	dma_cfg::gen2drv.put(tx);
	//wait for a clock in driver for data
	dma_cfg::drv2gen.get(rx);
	data = rx.data;
endtask : regs_read

// TODO : confirm prototype
// Write Register 
task regs_write(bit[3:0] address, bit [15:0] data);
	tx = new();
	tx.cs = 1'b0; 
	tx.ior = 1'b1;
	tx.iow = 1'b0;
	tx.addr_lo = address;
	tx.data = data;
	tx.dreq = 4'b0;
	tx.hlda = 1'b0; 
	tx.eop = 1'b1;
	tx.pkt_type = REG_WRITE;
	dma_cfg::gen2drv.put(tx);
endtask : regs_write
*/
// Constraints
	constraint dreq_c{
		dreq inside {[0:15]};
		dreq != dreq_old;
	}
	
	function void post_randomize();
		dreq_old = dreq;
	endfunction
	
// TODO: use rand variables for register fields
// TODO : Add constraints for other control signals
// Register Constraints
/*
constraint mode_reg_c {
	foreach(MODE_REG[i])  MODE_REG.mode_sel == 1;			// Only single  transfer mode supported
	foreach(MODE_REG[i])  MODE_REG.trans_type inside {1,2}; // Only read/write transfers supported
}

constraint cmd_reg_c {
	CMD_REG.mem2mem_en == 0;		// memory to memory transfers not supported
	CMD_REG.ch0_addr_hold == 0;		// Channel 0 address hold disabled
	CMD_REG.timing_type == 0; 		// Only normal timing_type supported
	CMD_REG.priority_type == 1; 	// Rotating priority_type supported
	CMD_REG.dreq_sense == 1;
	CMD_REG.dack_sense == 0;
}

constraint request_reg_c {
	REQ_REG.reserved == 0;
}

constraint mask_reg_c {
	MASK_REG.reserved == 0;
}
constraint transaction_c{
if(tx_type == REG_READ_CFG) {	cs = 1'b0; 
								ior = 1'b0;
								iow = 1'b1; 
								dreq = 4'b0;
								hlda = 1'b0;
								eop = 1'b1;}
else if(tx_type == REG_WRITE_CFG) 
							{	cs = 1'b0; 
								ior = 1'b1;
								iow = 1'b0;
								dreq = 4'b0;
								hlda = 1'b0;
								eop = 1'b1;}

}
*/
endclass : dma_transaction



// Order matters here so include in order of compilation dependencies

`include "dma_transaction.sv"
`include "dma_if.sv"
`include "dma_config.sv"
`include "dma_generator.sv"
`include "dma_driver.sv"
`include "dma_monitor.sv"
`include "dma_coverage.sv"
`include "dma_scoreboard.sv"
`include "dma_env.sv"
`include "dma_test.sv"
// `include "dma_assertions.sv"
`include "dma_datapath.sv"
`include "dma_priority.sv"
`include "dma_reg_file.sv"
`include "dma_control.sv"
`include "dma_reg_if.sv"
`include "dma_control_if.sv"
`include "dma_reg_pkg.sv"
`include "dma_top.sv"
`include "dma_tb_top.sv"
